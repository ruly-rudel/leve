
`define XLEN    64
`define FLEN    64
`define MXLEN   64
`define SXLEN   64
`define NUM_REG 32
`define FP_NUM_REG 32
`define NUM_CSR 4096
